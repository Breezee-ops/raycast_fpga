module sin(input [8:0] angle, output [9:0] val);



always_comb begin
case (angle)
9'd0 : val = 10'b0000100000;
9'd1 : val = 10'b0000011111;
9'd2 : val = 10'b0000011111;
9'd3 : val = 10'b0000011111;
9'd4 : val = 10'b0000011111;
9'd5 : val = 10'b0000011111;
9'd6 : val = 10'b0000011111;
9'd7 : val = 10'b0000011111;
9'd8 : val = 10'b0000011111;
9'd9 : val = 10'b0000011111;
9'd10 : val = 10'b0000011111;
9'd11 : val = 10'b0000011111;
9'd12 : val = 10'b0000011111;
9'd13 : val = 10'b0000011111;
9'd14 : val = 10'b0000011111;
9'd15 : val = 10'b0000011110;
9'd16 : val = 10'b0000011110;
9'd17 : val = 10'b0000011110;
9'd18 : val = 10'b0000011110;
9'd19 : val = 10'b0000011110;
9'd20 : val = 10'b0000011110;
9'd21 : val = 10'b0000011101;
9'd22 : val = 10'b0000011101;
9'd23 : val = 10'b0000011101;
9'd24 : val = 10'b0000011101;
9'd25 : val = 10'b0000011101;
9'd26 : val = 10'b0000011100;
9'd27 : val = 10'b0000011100;
9'd28 : val = 10'b0000011100;
9'd29 : val = 10'b0000011011;
9'd30 : val = 10'b0000011011;
9'd31 : val = 10'b0000011011;
9'd32 : val = 10'b0000011011;
9'd33 : val = 10'b0000011010;
9'd34 : val = 10'b0000011010;
9'd35 : val = 10'b0000011010;
9'd36 : val = 10'b0000011001;
9'd37 : val = 10'b0000011001;
9'd38 : val = 10'b0000011001;
9'd39 : val = 10'b0000011000;
9'd40 : val = 10'b0000011000;
9'd41 : val = 10'b0000011000;
9'd42 : val = 10'b0000010111;
9'd43 : val = 10'b0000010111;
9'd44 : val = 10'b0000010111;
9'd45 : val = 10'b0000010110;
9'd46 : val = 10'b0000010110;
9'd47 : val = 10'b0000010101;
9'd48 : val = 10'b0000010101;
9'd49 : val = 10'b0000010100;
9'd50 : val = 10'b0000010100;
9'd51 : val = 10'b0000010100;
9'd52 : val = 10'b0000010011;
9'd53 : val = 10'b0000010011;
9'd54 : val = 10'b0000010010;
9'd55 : val = 10'b0000010010;
9'd56 : val = 10'b0000010001;
9'd57 : val = 10'b0000010001;
9'd58 : val = 10'b0000010000;
9'd59 : val = 10'b0000010000;
9'd60 : val = 10'b0000010000;
9'd61 : val = 10'b0000001111;
9'd62 : val = 10'b0000001111;
9'd63 : val = 10'b0000001110;
9'd64 : val = 10'b0000001110;
9'd65 : val = 10'b0000001101;
9'd66 : val = 10'b0000001101;
9'd67 : val = 10'b0000001100;
9'd68 : val = 10'b0000001011;
9'd69 : val = 10'b0000001011;
9'd70 : val = 10'b0000001010;
9'd71 : val = 10'b0000001010;
9'd72 : val = 10'b0000001001;
9'd73 : val = 10'b0000001001;
9'd74 : val = 10'b0000001000;
9'd75 : val = 10'b0000001000;
9'd76 : val = 10'b0000000111;
9'd77 : val = 10'b0000000111;
9'd78 : val = 10'b0000000110;
9'd79 : val = 10'b0000000110;
9'd80 : val = 10'b0000000101;
9'd81 : val = 10'b0000000101;
9'd82 : val = 10'b0000000100;
9'd83 : val = 10'b0000000011;
9'd84 : val = 10'b0000000011;
9'd85 : val = 10'b0000000010;
9'd86 : val = 10'b0000000010;
9'd87 : val = 10'b0000000001;
9'd88 : val = 10'b0000000001;
9'd89 : val = 10'b0000000000;
9'd90 : val = 10'b0000000000;
9'd91 : val = 10'b0000000000;
9'd92 : val = 10'b1111111111;
9'd93 : val = 10'b1111111111;
9'd94 : val = 10'b1111111110;
9'd95 : val = 10'b1111111110;
9'd96 : val = 10'b1111111101;
9'd97 : val = 10'b1111111101;
9'd98 : val = 10'b1111111100;
9'd99 : val = 10'b1111111011;
9'd100 : val = 10'b1111111011;
9'd101 : val = 10'b1111111010;
9'd102 : val = 10'b1111111010;
9'd103 : val = 10'b1111111001;
9'd104 : val = 10'b1111111001;
9'd105 : val = 10'b1111111000;
9'd106 : val = 10'b1111111000;
9'd107 : val = 10'b1111110111;
9'd108 : val = 10'b1111110111;
9'd109 : val = 10'b1111110110;
9'd110 : val = 10'b1111110110;
9'd111 : val = 10'b1111110101;
9'd112 : val = 10'b1111110101;
9'd113 : val = 10'b1111110100;
9'd114 : val = 10'b1111110011;
9'd115 : val = 10'b1111110011;
9'd116 : val = 10'b1111110010;
9'd117 : val = 10'b1111110010;
9'd118 : val = 10'b1111110001;
9'd119 : val = 10'b1111110001;
9'd120 : val = 10'b1111110001;
9'd121 : val = 10'b1111110000;
9'd122 : val = 10'b1111110000;
9'd123 : val = 10'b1111101111;
9'd124 : val = 10'b1111101111;
9'd125 : val = 10'b1111101110;
9'd126 : val = 10'b1111101110;
9'd127 : val = 10'b1111101101;
9'd128 : val = 10'b1111101101;
9'd129 : val = 10'b1111101100;
9'd130 : val = 10'b1111101100;
9'd131 : val = 10'b1111101100;
9'd132 : val = 10'b1111101011;
9'd133 : val = 10'b1111101011;
9'd134 : val = 10'b1111101010;
9'd135 : val = 10'b1111101010;
9'd136 : val = 10'b1111101001;
9'd137 : val = 10'b1111101001;
9'd138 : val = 10'b1111101001;
9'd139 : val = 10'b1111101000;
9'd140 : val = 10'b1111101000;
9'd141 : val = 10'b1111101000;
9'd142 : val = 10'b1111100111;
9'd143 : val = 10'b1111100111;
9'd144 : val = 10'b1111100111;
9'd145 : val = 10'b1111100110;
9'd146 : val = 10'b1111100110;
9'd147 : val = 10'b1111100110;
9'd148 : val = 10'b1111100101;
9'd149 : val = 10'b1111100101;
9'd150 : val = 10'b1111100101;
9'd151 : val = 10'b1111100101;
9'd152 : val = 10'b1111100100;
9'd153 : val = 10'b1111100100;
9'd154 : val = 10'b1111100100;
9'd155 : val = 10'b1111100011;
9'd156 : val = 10'b1111100011;
9'd157 : val = 10'b1111100011;
9'd158 : val = 10'b1111100011;
9'd159 : val = 10'b1111100011;
9'd160 : val = 10'b1111100010;
9'd161 : val = 10'b1111100010;
9'd162 : val = 10'b1111100010;
9'd163 : val = 10'b1111100010;
9'd164 : val = 10'b1111100010;
9'd165 : val = 10'b1111100010;
9'd166 : val = 10'b1111100001;
9'd167 : val = 10'b1111100001;
9'd168 : val = 10'b1111100001;
9'd169 : val = 10'b1111100001;
9'd170 : val = 10'b1111100001;
9'd171 : val = 10'b1111100001;
9'd172 : val = 10'b1111100001;
9'd173 : val = 10'b1111100001;
9'd174 : val = 10'b1111100001;
9'd175 : val = 10'b1111100001;
9'd176 : val = 10'b1111100001;
9'd177 : val = 10'b1111100001;
9'd178 : val = 10'b1111100001;
9'd179 : val = 10'b1111100001;
9'd180 : val = 10'b1111100000;
9'd181 : val = 10'b1111100001;
9'd182 : val = 10'b1111100001;
9'd183 : val = 10'b1111100001;
9'd184 : val = 10'b1111100001;
9'd185 : val = 10'b1111100001;
9'd186 : val = 10'b1111100001;
9'd187 : val = 10'b1111100001;
9'd188 : val = 10'b1111100001;
9'd189 : val = 10'b1111100001;
9'd190 : val = 10'b1111100001;
9'd191 : val = 10'b1111100001;
9'd192 : val = 10'b1111100001;
9'd193 : val = 10'b1111100001;
9'd194 : val = 10'b1111100001;
9'd195 : val = 10'b1111100010;
9'd196 : val = 10'b1111100010;
9'd197 : val = 10'b1111100010;
9'd198 : val = 10'b1111100010;
9'd199 : val = 10'b1111100010;
9'd200 : val = 10'b1111100010;
9'd201 : val = 10'b1111100011;
9'd202 : val = 10'b1111100011;
9'd203 : val = 10'b1111100011;
9'd204 : val = 10'b1111100011;
9'd205 : val = 10'b1111100011;
9'd206 : val = 10'b1111100100;
9'd207 : val = 10'b1111100100;
9'd208 : val = 10'b1111100100;
9'd209 : val = 10'b1111100101;
9'd210 : val = 10'b1111100101;
9'd211 : val = 10'b1111100101;
9'd212 : val = 10'b1111100101;
9'd213 : val = 10'b1111100110;
9'd214 : val = 10'b1111100110;
9'd215 : val = 10'b1111100110;
9'd216 : val = 10'b1111100111;
9'd217 : val = 10'b1111100111;
9'd218 : val = 10'b1111100111;
9'd219 : val = 10'b1111101000;
9'd220 : val = 10'b1111101000;
9'd221 : val = 10'b1111101000;
9'd222 : val = 10'b1111101001;
9'd223 : val = 10'b1111101001;
9'd224 : val = 10'b1111101001;
9'd225 : val = 10'b1111101010;
9'd226 : val = 10'b1111101010;
9'd227 : val = 10'b1111101011;
9'd228 : val = 10'b1111101011;
9'd229 : val = 10'b1111101100;
9'd230 : val = 10'b1111101100;
9'd231 : val = 10'b1111101100;
9'd232 : val = 10'b1111101101;
9'd233 : val = 10'b1111101101;
9'd234 : val = 10'b1111101110;
9'd235 : val = 10'b1111101110;
9'd236 : val = 10'b1111101111;
9'd237 : val = 10'b1111101111;
9'd238 : val = 10'b1111110000;
9'd239 : val = 10'b1111110000;
9'd240 : val = 10'b1111110000;
9'd241 : val = 10'b1111110001;
9'd242 : val = 10'b1111110001;
9'd243 : val = 10'b1111110010;
9'd244 : val = 10'b1111110010;
9'd245 : val = 10'b1111110011;
9'd246 : val = 10'b1111110011;
9'd247 : val = 10'b1111110100;
9'd248 : val = 10'b1111110101;
9'd249 : val = 10'b1111110101;
9'd250 : val = 10'b1111110110;
9'd251 : val = 10'b1111110110;
9'd252 : val = 10'b1111110111;
9'd253 : val = 10'b1111110111;
9'd254 : val = 10'b1111111000;
9'd255 : val = 10'b1111111000;
9'd256 : val = 10'b1111111001;
9'd257 : val = 10'b1111111001;
9'd258 : val = 10'b1111111010;
9'd259 : val = 10'b1111111010;
9'd260 : val = 10'b1111111011;
9'd261 : val = 10'b1111111011;
9'd262 : val = 10'b1111111100;
9'd263 : val = 10'b1111111101;
9'd264 : val = 10'b1111111101;
9'd265 : val = 10'b1111111110;
9'd266 : val = 10'b1111111110;
9'd267 : val = 10'b1111111111;
9'd268 : val = 10'b1111111111;
9'd269 : val = 10'b0000000000;
9'd270 : val = 10'b0000000000;
9'd271 : val = 10'b0000000000;
9'd272 : val = 10'b0000000001;
9'd273 : val = 10'b0000000001;
9'd274 : val = 10'b0000000010;
9'd275 : val = 10'b0000000010;
9'd276 : val = 10'b0000000011;
9'd277 : val = 10'b0000000011;
9'd278 : val = 10'b0000000100;
9'd279 : val = 10'b0000000101;
9'd280 : val = 10'b0000000101;
9'd281 : val = 10'b0000000110;
9'd282 : val = 10'b0000000110;
9'd283 : val = 10'b0000000111;
9'd284 : val = 10'b0000000111;
9'd285 : val = 10'b0000001000;
9'd286 : val = 10'b0000001000;
9'd287 : val = 10'b0000001001;
9'd288 : val = 10'b0000001001;
9'd289 : val = 10'b0000001010;
9'd290 : val = 10'b0000001010;
9'd291 : val = 10'b0000001011;
9'd292 : val = 10'b0000001011;
9'd293 : val = 10'b0000001100;
9'd294 : val = 10'b0000001101;
9'd295 : val = 10'b0000001101;
9'd296 : val = 10'b0000001110;
9'd297 : val = 10'b0000001110;
9'd298 : val = 10'b0000001111;
9'd299 : val = 10'b0000001111;
9'd300 : val = 10'b0000010000;
9'd301 : val = 10'b0000010000;
9'd302 : val = 10'b0000010000;
9'd303 : val = 10'b0000010001;
9'd304 : val = 10'b0000010001;
9'd305 : val = 10'b0000010010;
9'd306 : val = 10'b0000010010;
9'd307 : val = 10'b0000010011;
9'd308 : val = 10'b0000010011;
9'd309 : val = 10'b0000010100;
9'd310 : val = 10'b0000010100;
9'd311 : val = 10'b0000010100;
9'd312 : val = 10'b0000010101;
9'd313 : val = 10'b0000010101;
9'd314 : val = 10'b0000010110;
9'd315 : val = 10'b0000010110;
9'd316 : val = 10'b0000010111;
9'd317 : val = 10'b0000010111;
9'd318 : val = 10'b0000010111;
9'd319 : val = 10'b0000011000;
9'd320 : val = 10'b0000011000;
9'd321 : val = 10'b0000011000;
9'd322 : val = 10'b0000011001;
9'd323 : val = 10'b0000011001;
9'd324 : val = 10'b0000011001;
9'd325 : val = 10'b0000011010;
9'd326 : val = 10'b0000011010;
9'd327 : val = 10'b0000011010;
9'd328 : val = 10'b0000011011;
9'd329 : val = 10'b0000011011;
9'd330 : val = 10'b0000011011;
9'd331 : val = 10'b0000011011;
9'd332 : val = 10'b0000011100;
9'd333 : val = 10'b0000011100;
9'd334 : val = 10'b0000011100;
9'd335 : val = 10'b0000011101;
9'd336 : val = 10'b0000011101;
9'd337 : val = 10'b0000011101;
9'd338 : val = 10'b0000011101;
9'd339 : val = 10'b0000011101;
9'd340 : val = 10'b0000011110;
9'd341 : val = 10'b0000011110;
9'd342 : val = 10'b0000011110;
9'd343 : val = 10'b0000011110;
9'd344 : val = 10'b0000011110;
9'd345 : val = 10'b0000011110;
9'd346 : val = 10'b0000011111;
9'd347 : val = 10'b0000011111;
9'd348 : val = 10'b0000011111;
9'd349 : val = 10'b0000011111;
9'd350 : val = 10'b0000011111;
9'd351 : val = 10'b0000011111;
9'd352 : val = 10'b0000011111;
9'd353 : val = 10'b0000011111;
9'd354 : val = 10'b0000011111;
9'd355 : val = 10'b0000011111;
9'd356 : val = 10'b0000011111;
9'd357 : val = 10'b0000011111;
9'd358 : val = 10'b0000011111;
9'd359 : val = 10'b0000011111;
default: val = 10'd0;
endcase
end
endmodule
